// testbench for fulladder using oop
-------------‐-----------
-------------‐-----------
class 